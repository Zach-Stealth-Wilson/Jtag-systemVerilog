/*
 * Copyright (c) 2024 Your Name
 * SPDX-License-Identifier: Apache-2.0
 */

`default_nettype none

module tt_um_example (
    input  wire [7:0] ui_in,    // Dedicated inputs
    output wire [7:0] uo_out,   // Dedicated outputs
    input  wire [7:0] uio_in,   // IOs: Input path
    output wire [7:0] uio_out,  // IOs: Output path
    output wire [7:0] uio_oe,   // IOs: Enable path (active high: 0=input, 1=output)
    input  wire       ena,      // always 1 when the design is powered, so you can ignore it
    input  wire       clk,      // clock
    input  wire       rst_n     // reset_n - low to reset
);

  // All output pins must be assigned. If not used, assign to 0.
  
  assign uio_out = 0;
  assign uio_oe  = 0;

  // List all unused inputs to prevent warnings .a(ui_in[7:0]), .b(uio_in[7:0])
  wire _unused = &{ena, clk, rst_n, 1'b0};

    tt_um_jtag_test_logic top(.tck(clk), .tms(), .tdi(), .reset(rst_n), .tdo(uo_out[0]), .bsr_tdi(), .bsr_clk(), .bsr_update(), .bsr_shift(), .bsr_mode(), .bsr_tdo(), .sys_clk(), .dbg_clk(), .dm_reset() );

endmodule
